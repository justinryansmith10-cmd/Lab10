module seven_segment_negative(i,o);

input i;
output reg [6:0]o; 

// HEX out - rewire DE1
//  ---0---
// |       |
// 5       1
// |       |
//  ---6---
// |       |
// 4       2
// |       |
//  ---3---

endmodule